module decoder(
	input wire[31:0] inst,
	input wire reset,					// Pone todas las salidas en 0
	output wire[4:0] rd,
	output wire[4:0] rs1,
	output wire[4:0] rs2,
	output wire[2:0] funct3,
	output reg rd_enc,				// Habilita que el valor del bus C se guarde en el registro rd
	output reg rs1_ena,				// Habilita que el valor del registro rs1 se copie al bus A
	output reg rs2_enb,				// Habilita que el valor del registro rs2 se copie al bus B
	output reg imm_en,				// Habilita el calculo de imm y su copia al bus IMM
	output reg imm_enb,				// Habilita que el valor del imm se copie al bus B
	//output wire pc_ena,
	output reg ALU_en,				// Habilita la ALU
	output wire ALU_flag,			// Flag para ciertas operaciones de la ALU
	output reg mem_en,				// Habilita el acceso a memoria
	output wire rw,					// Indica si el acceso a memoria es de lectura o escritura
	output reg is_jmp,
	output reg is_fence,
	output reg is_system,
	output reg is_invalid
);


wire[4:0] opcode = reset ? 5'b11111 : inst[6:2];
assign rd = inst[11:7];
assign funct3 = inst[14:12];
assign rs1 = inst[19:15];
assign rs2 = inst[24:20];
assign ALU_flag = inst[30];
assign rw = inst[5];				// rw = 1 si es STORE, = 0 si es LOAD

always @(opcode)
begin
    case(opcode)
		  // LUI (U) o AIUPC(U)
        5'b01101, 5'b00101: begin
			  ALU_en = 1'b1;
			  rd_enc = 1'b1;				  
			  //rs1 = (opcode[3] == 1'b1) ? 5'b00000 : rs1;	// ???? Puedo redefinir rs1 así? rd = 0 + imm si es LUI
			  rs1_ena = opcode[3];
			  // PC_ena = !opcode[3];	// Mandar el PC al A si es AIUPC ?
			  imm_en = 1'b1;
			  imm_enb = 1'b1;
			  rs2_enb = 1'b0;
			  mem_en = 1'b0;
			  is_jmp = 1'b0;
			  is_fence = 1'b0;
			  is_system = 1'b0;
			  is_invalid = 1'b0;
			end
		  // JAL (J), JALR (I) o BRANCH (B)
		  5'b11011, 5'b11001, 5'b11000: begin		
			  is_jmp = 1'b1;
			  imm_en = 1'b1;				// !!!! El imm no debería ir a la ALU sino al Jmp Ctrl
			  rs1_ena = !opcode[1];		// !!!! El rs1 debería ir al Jmp Ctrl ya que add = rs1 + imm en JALR y BRANCH
			  ALU_en = !opcode[0];		// ALU_en = 1 si es BRANCH
			  //rs1_ena = !opcode[0];	// !!!! Pero si es BRANCH rs1 también tiene que ir a la ALU
			  rs2_enb = !opcode[0];		// rs2_enb = 1 si es BRANCH
			  // TODO: Chequear funct3
			  rd_enc = 1'b0;
			  imm_enb = 1'b0;
			  mem_en = 1'b0;
			  is_fence = 1'b0;
			  is_system = 1'b0;
			  is_invalid = 1'b0;
		  end
		  //  LOAD (I) o STORE (S)
		  5'b00000, 5'b01000: begin	
			  mem_en = 1'b1;
			  rs1_ena = 1'b1;				// !!!! El rs1 debería ir al Address Builder ya que add = rs1 + imm en LOAD y STORE
			  imm_en = 1'b1;				// !!!! El imm debería ir al Address Builder
			  rs2_enb = opcode[3];		// !!!! El rs2 debería ir al Memory Manager(? si es STORE
			  rd_enc = !opcode[3];		// rd_enc = 1 si es LOAD
			  imm_enb = 1'b0;
			  ALU_en = 1'b0;
			  is_jmp = 1'b0;
			  is_fence = 1'b0;
			  is_system = 1'b0;
			  is_invalid = 1'b0;
		  end
		  // ALUI (I) o ALU (R)
		  5'b00100, 5'b01100: begin
			  ALU_en = 1'b1;
			  rd_enc = 1'b1;
			  rs1_ena = 1'b1;
			  rs2_enb = opcode[3];		// rs2_enb = 1 si es ALU, = 0 si es ALUI
			  imm_en = !opcode[3];
			  imm_enb = !opcode[3];		// imm_enb = 1 si es ALUI, = 0 si es ALU
			  mem_en = 1'b0;
			  is_jmp = 1'b0;
			  is_fence = 1'b0;
			  is_system = 1'b0;
			  is_invalid = 1'b0;
		  end
		  // FENCE (R) or SYSTEM (R)
		  5'b00011, 5'b11100: begin		
			  is_fence = opcode[0];	
			  is_system = opcode[4];
			  rd_enc = 1'b0;
			  rs1_ena = 1'b0;
			  rs2_enb = 1'b0;
			  imm_en = 1'b0;
			  imm_enb = 1'b0;
			  ALU_en = 1'b0;
			  mem_en = 1'b0;
			  is_jmp = 1'b0;
			  is_invalid = 1'b0;
		  end
        default: begin 	// Invalid opcode
			  is_invalid = 1'b1;
			  rd_enc = 1'b0;
			  rs1_ena = 1'b0;
			  rs2_enb = 1'b0;
			  imm_en = 1'b0;
			  imm_enb = 1'b0;
			  ALU_en = 1'b0;
			  mem_en = 1'b0;
			  is_jmp = 1'b0;
			  is_fence = 1'b0;
			  is_system = 1'b0;
		  end
    endcase
end

endmodule