// megafunction wizard: %LPM_DECODE%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_DECODE 

// ============================================================
// File Name: peripheral_addr_dec.v
// Megafunction Name(s):
// 			LPM_DECODE
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 23.1std.0 Build 991 11/28/2023 SC Lite Edition
// ************************************************************

//Copyright (C) 2023  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and any partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details, at
//https://fpgasoftware.intel.com/eula.

module peripheral_addr_dec (
	data,
	enable,
	eq0,
	eq1,
	eq10,
	eq11,
	eq12,
	eq13,
	eq14,
	eq15,
	eq16,
	eq17,
	eq18,
	eq19,
	eq2,
	eq20,
	eq21,
	eq22,
	eq23,
	eq24,
	eq25,
	eq26,
	eq27,
	eq28,
	eq29,
	eq3,
	eq30,
	eq31,
	eq32,
	eq33,
	eq34,
	eq35,
	eq36,
	eq37,
	eq38,
	eq39,
	eq4,
	eq40,
	eq41,
	eq42,
	eq43,
	eq44,
	eq45,
	eq46,
	eq47,
	eq48,
	eq49,
	eq5,
	eq50,
	eq51,
	eq52,
	eq53,
	eq54,
	eq55,
	eq56,
	eq57,
	eq58,
	eq59,
	eq6,
	eq60,
	eq61,
	eq62,
	eq63,
	eq7,
	eq8,
	eq9);

	input	[5:0]  data;
	input	  enable;
	output	  eq0;
	output	  eq1;
	output	  eq10;
	output	  eq11;
	output	  eq12;
	output	  eq13;
	output	  eq14;
	output	  eq15;
	output	  eq16;
	output	  eq17;
	output	  eq18;
	output	  eq19;
	output	  eq2;
	output	  eq20;
	output	  eq21;
	output	  eq22;
	output	  eq23;
	output	  eq24;
	output	  eq25;
	output	  eq26;
	output	  eq27;
	output	  eq28;
	output	  eq29;
	output	  eq3;
	output	  eq30;
	output	  eq31;
	output	  eq32;
	output	  eq33;
	output	  eq34;
	output	  eq35;
	output	  eq36;
	output	  eq37;
	output	  eq38;
	output	  eq39;
	output	  eq4;
	output	  eq40;
	output	  eq41;
	output	  eq42;
	output	  eq43;
	output	  eq44;
	output	  eq45;
	output	  eq46;
	output	  eq47;
	output	  eq48;
	output	  eq49;
	output	  eq5;
	output	  eq50;
	output	  eq51;
	output	  eq52;
	output	  eq53;
	output	  eq54;
	output	  eq55;
	output	  eq56;
	output	  eq57;
	output	  eq58;
	output	  eq59;
	output	  eq6;
	output	  eq60;
	output	  eq61;
	output	  eq62;
	output	  eq63;
	output	  eq7;
	output	  eq8;
	output	  eq9;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: BaseDec NUMERIC "1"
// Retrieval info: PRIVATE: EnableInput NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "0"
// Retrieval info: PRIVATE: Latency NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: aclr NUMERIC "0"
// Retrieval info: PRIVATE: clken NUMERIC "0"
// Retrieval info: PRIVATE: eq0 NUMERIC "1"
// Retrieval info: PRIVATE: eq1 NUMERIC "1"
// Retrieval info: PRIVATE: eq10 NUMERIC "1"
// Retrieval info: PRIVATE: eq11 NUMERIC "1"
// Retrieval info: PRIVATE: eq12 NUMERIC "1"
// Retrieval info: PRIVATE: eq13 NUMERIC "1"
// Retrieval info: PRIVATE: eq14 NUMERIC "1"
// Retrieval info: PRIVATE: eq15 NUMERIC "1"
// Retrieval info: PRIVATE: eq16 NUMERIC "1"
// Retrieval info: PRIVATE: eq17 NUMERIC "1"
// Retrieval info: PRIVATE: eq18 NUMERIC "1"
// Retrieval info: PRIVATE: eq19 NUMERIC "1"
// Retrieval info: PRIVATE: eq2 NUMERIC "1"
// Retrieval info: PRIVATE: eq20 NUMERIC "1"
// Retrieval info: PRIVATE: eq21 NUMERIC "1"
// Retrieval info: PRIVATE: eq22 NUMERIC "1"
// Retrieval info: PRIVATE: eq23 NUMERIC "1"
// Retrieval info: PRIVATE: eq24 NUMERIC "1"
// Retrieval info: PRIVATE: eq25 NUMERIC "1"
// Retrieval info: PRIVATE: eq26 NUMERIC "1"
// Retrieval info: PRIVATE: eq27 NUMERIC "1"
// Retrieval info: PRIVATE: eq28 NUMERIC "1"
// Retrieval info: PRIVATE: eq29 NUMERIC "1"
// Retrieval info: PRIVATE: eq3 NUMERIC "1"
// Retrieval info: PRIVATE: eq30 NUMERIC "1"
// Retrieval info: PRIVATE: eq31 NUMERIC "1"
// Retrieval info: PRIVATE: eq32 NUMERIC "1"
// Retrieval info: PRIVATE: eq33 NUMERIC "1"
// Retrieval info: PRIVATE: eq34 NUMERIC "1"
// Retrieval info: PRIVATE: eq35 NUMERIC "1"
// Retrieval info: PRIVATE: eq36 NUMERIC "1"
// Retrieval info: PRIVATE: eq37 NUMERIC "1"
// Retrieval info: PRIVATE: eq38 NUMERIC "1"
// Retrieval info: PRIVATE: eq39 NUMERIC "1"
// Retrieval info: PRIVATE: eq4 NUMERIC "1"
// Retrieval info: PRIVATE: eq40 NUMERIC "1"
// Retrieval info: PRIVATE: eq41 NUMERIC "1"
// Retrieval info: PRIVATE: eq42 NUMERIC "1"
// Retrieval info: PRIVATE: eq43 NUMERIC "1"
// Retrieval info: PRIVATE: eq44 NUMERIC "1"
// Retrieval info: PRIVATE: eq45 NUMERIC "1"
// Retrieval info: PRIVATE: eq46 NUMERIC "1"
// Retrieval info: PRIVATE: eq47 NUMERIC "1"
// Retrieval info: PRIVATE: eq48 NUMERIC "1"
// Retrieval info: PRIVATE: eq49 NUMERIC "1"
// Retrieval info: PRIVATE: eq5 NUMERIC "1"
// Retrieval info: PRIVATE: eq50 NUMERIC "1"
// Retrieval info: PRIVATE: eq51 NUMERIC "1"
// Retrieval info: PRIVATE: eq52 NUMERIC "1"
// Retrieval info: PRIVATE: eq53 NUMERIC "1"
// Retrieval info: PRIVATE: eq54 NUMERIC "1"
// Retrieval info: PRIVATE: eq55 NUMERIC "1"
// Retrieval info: PRIVATE: eq56 NUMERIC "1"
// Retrieval info: PRIVATE: eq57 NUMERIC "1"
// Retrieval info: PRIVATE: eq58 NUMERIC "1"
// Retrieval info: PRIVATE: eq59 NUMERIC "1"
// Retrieval info: PRIVATE: eq6 NUMERIC "1"
// Retrieval info: PRIVATE: eq60 NUMERIC "1"
// Retrieval info: PRIVATE: eq61 NUMERIC "1"
// Retrieval info: PRIVATE: eq62 NUMERIC "1"
// Retrieval info: PRIVATE: eq63 NUMERIC "1"
// Retrieval info: PRIVATE: eq7 NUMERIC "1"
// Retrieval info: PRIVATE: eq8 NUMERIC "1"
// Retrieval info: PRIVATE: eq9 NUMERIC "1"
// Retrieval info: PRIVATE: nBit NUMERIC "6"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_DECODES NUMERIC "64"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DECODE"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "6"
// Retrieval info: USED_PORT: @eq 0 0 64 0 OUTPUT NODEFVAL "@eq[63..0]"
// Retrieval info: USED_PORT: data 0 0 6 0 INPUT NODEFVAL "data[5..0]"
// Retrieval info: USED_PORT: enable 0 0 0 0 INPUT NODEFVAL "enable"
// Retrieval info: USED_PORT: eq0 0 0 0 0 OUTPUT NODEFVAL "eq0"
// Retrieval info: USED_PORT: eq1 0 0 0 0 OUTPUT NODEFVAL "eq1"
// Retrieval info: USED_PORT: eq10 0 0 0 0 OUTPUT NODEFVAL "eq10"
// Retrieval info: USED_PORT: eq11 0 0 0 0 OUTPUT NODEFVAL "eq11"
// Retrieval info: USED_PORT: eq12 0 0 0 0 OUTPUT NODEFVAL "eq12"
// Retrieval info: USED_PORT: eq13 0 0 0 0 OUTPUT NODEFVAL "eq13"
// Retrieval info: USED_PORT: eq14 0 0 0 0 OUTPUT NODEFVAL "eq14"
// Retrieval info: USED_PORT: eq15 0 0 0 0 OUTPUT NODEFVAL "eq15"
// Retrieval info: USED_PORT: eq16 0 0 0 0 OUTPUT NODEFVAL "eq16"
// Retrieval info: USED_PORT: eq17 0 0 0 0 OUTPUT NODEFVAL "eq17"
// Retrieval info: USED_PORT: eq18 0 0 0 0 OUTPUT NODEFVAL "eq18"
// Retrieval info: USED_PORT: eq19 0 0 0 0 OUTPUT NODEFVAL "eq19"
// Retrieval info: USED_PORT: eq2 0 0 0 0 OUTPUT NODEFVAL "eq2"
// Retrieval info: USED_PORT: eq20 0 0 0 0 OUTPUT NODEFVAL "eq20"
// Retrieval info: USED_PORT: eq21 0 0 0 0 OUTPUT NODEFVAL "eq21"
// Retrieval info: USED_PORT: eq22 0 0 0 0 OUTPUT NODEFVAL "eq22"
// Retrieval info: USED_PORT: eq23 0 0 0 0 OUTPUT NODEFVAL "eq23"
// Retrieval info: USED_PORT: eq24 0 0 0 0 OUTPUT NODEFVAL "eq24"
// Retrieval info: USED_PORT: eq25 0 0 0 0 OUTPUT NODEFVAL "eq25"
// Retrieval info: USED_PORT: eq26 0 0 0 0 OUTPUT NODEFVAL "eq26"
// Retrieval info: USED_PORT: eq27 0 0 0 0 OUTPUT NODEFVAL "eq27"
// Retrieval info: USED_PORT: eq28 0 0 0 0 OUTPUT NODEFVAL "eq28"
// Retrieval info: USED_PORT: eq29 0 0 0 0 OUTPUT NODEFVAL "eq29"
// Retrieval info: USED_PORT: eq3 0 0 0 0 OUTPUT NODEFVAL "eq3"
// Retrieval info: USED_PORT: eq30 0 0 0 0 OUTPUT NODEFVAL "eq30"
// Retrieval info: USED_PORT: eq31 0 0 0 0 OUTPUT NODEFVAL "eq31"
// Retrieval info: USED_PORT: eq32 0 0 0 0 OUTPUT NODEFVAL "eq32"
// Retrieval info: USED_PORT: eq33 0 0 0 0 OUTPUT NODEFVAL "eq33"
// Retrieval info: USED_PORT: eq34 0 0 0 0 OUTPUT NODEFVAL "eq34"
// Retrieval info: USED_PORT: eq35 0 0 0 0 OUTPUT NODEFVAL "eq35"
// Retrieval info: USED_PORT: eq36 0 0 0 0 OUTPUT NODEFVAL "eq36"
// Retrieval info: USED_PORT: eq37 0 0 0 0 OUTPUT NODEFVAL "eq37"
// Retrieval info: USED_PORT: eq38 0 0 0 0 OUTPUT NODEFVAL "eq38"
// Retrieval info: USED_PORT: eq39 0 0 0 0 OUTPUT NODEFVAL "eq39"
// Retrieval info: USED_PORT: eq4 0 0 0 0 OUTPUT NODEFVAL "eq4"
// Retrieval info: USED_PORT: eq40 0 0 0 0 OUTPUT NODEFVAL "eq40"
// Retrieval info: USED_PORT: eq41 0 0 0 0 OUTPUT NODEFVAL "eq41"
// Retrieval info: USED_PORT: eq42 0 0 0 0 OUTPUT NODEFVAL "eq42"
// Retrieval info: USED_PORT: eq43 0 0 0 0 OUTPUT NODEFVAL "eq43"
// Retrieval info: USED_PORT: eq44 0 0 0 0 OUTPUT NODEFVAL "eq44"
// Retrieval info: USED_PORT: eq45 0 0 0 0 OUTPUT NODEFVAL "eq45"
// Retrieval info: USED_PORT: eq46 0 0 0 0 OUTPUT NODEFVAL "eq46"
// Retrieval info: USED_PORT: eq47 0 0 0 0 OUTPUT NODEFVAL "eq47"
// Retrieval info: USED_PORT: eq48 0 0 0 0 OUTPUT NODEFVAL "eq48"
// Retrieval info: USED_PORT: eq49 0 0 0 0 OUTPUT NODEFVAL "eq49"
// Retrieval info: USED_PORT: eq5 0 0 0 0 OUTPUT NODEFVAL "eq5"
// Retrieval info: USED_PORT: eq50 0 0 0 0 OUTPUT NODEFVAL "eq50"
// Retrieval info: USED_PORT: eq51 0 0 0 0 OUTPUT NODEFVAL "eq51"
// Retrieval info: USED_PORT: eq52 0 0 0 0 OUTPUT NODEFVAL "eq52"
// Retrieval info: USED_PORT: eq53 0 0 0 0 OUTPUT NODEFVAL "eq53"
// Retrieval info: USED_PORT: eq54 0 0 0 0 OUTPUT NODEFVAL "eq54"
// Retrieval info: USED_PORT: eq55 0 0 0 0 OUTPUT NODEFVAL "eq55"
// Retrieval info: USED_PORT: eq56 0 0 0 0 OUTPUT NODEFVAL "eq56"
// Retrieval info: USED_PORT: eq57 0 0 0 0 OUTPUT NODEFVAL "eq57"
// Retrieval info: USED_PORT: eq58 0 0 0 0 OUTPUT NODEFVAL "eq58"
// Retrieval info: USED_PORT: eq59 0 0 0 0 OUTPUT NODEFVAL "eq59"
// Retrieval info: USED_PORT: eq6 0 0 0 0 OUTPUT NODEFVAL "eq6"
// Retrieval info: USED_PORT: eq60 0 0 0 0 OUTPUT NODEFVAL "eq60"
// Retrieval info: USED_PORT: eq61 0 0 0 0 OUTPUT NODEFVAL "eq61"
// Retrieval info: USED_PORT: eq62 0 0 0 0 OUTPUT NODEFVAL "eq62"
// Retrieval info: USED_PORT: eq63 0 0 0 0 OUTPUT NODEFVAL "eq63"
// Retrieval info: USED_PORT: eq7 0 0 0 0 OUTPUT NODEFVAL "eq7"
// Retrieval info: USED_PORT: eq8 0 0 0 0 OUTPUT NODEFVAL "eq8"
// Retrieval info: USED_PORT: eq9 0 0 0 0 OUTPUT NODEFVAL "eq9"
// Retrieval info: CONNECT: @data 0 0 6 0 data 0 0 6 0
// Retrieval info: CONNECT: @enable 0 0 0 0 enable 0 0 0 0
// Retrieval info: CONNECT: eq0 0 0 0 0 @eq 0 0 1 0
// Retrieval info: CONNECT: eq1 0 0 0 0 @eq 0 0 1 1
// Retrieval info: CONNECT: eq10 0 0 0 0 @eq 0 0 1 10
// Retrieval info: CONNECT: eq11 0 0 0 0 @eq 0 0 1 11
// Retrieval info: CONNECT: eq12 0 0 0 0 @eq 0 0 1 12
// Retrieval info: CONNECT: eq13 0 0 0 0 @eq 0 0 1 13
// Retrieval info: CONNECT: eq14 0 0 0 0 @eq 0 0 1 14
// Retrieval info: CONNECT: eq15 0 0 0 0 @eq 0 0 1 15
// Retrieval info: CONNECT: eq16 0 0 0 0 @eq 0 0 1 16
// Retrieval info: CONNECT: eq17 0 0 0 0 @eq 0 0 1 17
// Retrieval info: CONNECT: eq18 0 0 0 0 @eq 0 0 1 18
// Retrieval info: CONNECT: eq19 0 0 0 0 @eq 0 0 1 19
// Retrieval info: CONNECT: eq2 0 0 0 0 @eq 0 0 1 2
// Retrieval info: CONNECT: eq20 0 0 0 0 @eq 0 0 1 20
// Retrieval info: CONNECT: eq21 0 0 0 0 @eq 0 0 1 21
// Retrieval info: CONNECT: eq22 0 0 0 0 @eq 0 0 1 22
// Retrieval info: CONNECT: eq23 0 0 0 0 @eq 0 0 1 23
// Retrieval info: CONNECT: eq24 0 0 0 0 @eq 0 0 1 24
// Retrieval info: CONNECT: eq25 0 0 0 0 @eq 0 0 1 25
// Retrieval info: CONNECT: eq26 0 0 0 0 @eq 0 0 1 26
// Retrieval info: CONNECT: eq27 0 0 0 0 @eq 0 0 1 27
// Retrieval info: CONNECT: eq28 0 0 0 0 @eq 0 0 1 28
// Retrieval info: CONNECT: eq29 0 0 0 0 @eq 0 0 1 29
// Retrieval info: CONNECT: eq3 0 0 0 0 @eq 0 0 1 3
// Retrieval info: CONNECT: eq30 0 0 0 0 @eq 0 0 1 30
// Retrieval info: CONNECT: eq31 0 0 0 0 @eq 0 0 1 31
// Retrieval info: CONNECT: eq32 0 0 0 0 @eq 0 0 1 32
// Retrieval info: CONNECT: eq33 0 0 0 0 @eq 0 0 1 33
// Retrieval info: CONNECT: eq34 0 0 0 0 @eq 0 0 1 34
// Retrieval info: CONNECT: eq35 0 0 0 0 @eq 0 0 1 35
// Retrieval info: CONNECT: eq36 0 0 0 0 @eq 0 0 1 36
// Retrieval info: CONNECT: eq37 0 0 0 0 @eq 0 0 1 37
// Retrieval info: CONNECT: eq38 0 0 0 0 @eq 0 0 1 38
// Retrieval info: CONNECT: eq39 0 0 0 0 @eq 0 0 1 39
// Retrieval info: CONNECT: eq4 0 0 0 0 @eq 0 0 1 4
// Retrieval info: CONNECT: eq40 0 0 0 0 @eq 0 0 1 40
// Retrieval info: CONNECT: eq41 0 0 0 0 @eq 0 0 1 41
// Retrieval info: CONNECT: eq42 0 0 0 0 @eq 0 0 1 42
// Retrieval info: CONNECT: eq43 0 0 0 0 @eq 0 0 1 43
// Retrieval info: CONNECT: eq44 0 0 0 0 @eq 0 0 1 44
// Retrieval info: CONNECT: eq45 0 0 0 0 @eq 0 0 1 45
// Retrieval info: CONNECT: eq46 0 0 0 0 @eq 0 0 1 46
// Retrieval info: CONNECT: eq47 0 0 0 0 @eq 0 0 1 47
// Retrieval info: CONNECT: eq48 0 0 0 0 @eq 0 0 1 48
// Retrieval info: CONNECT: eq49 0 0 0 0 @eq 0 0 1 49
// Retrieval info: CONNECT: eq5 0 0 0 0 @eq 0 0 1 5
// Retrieval info: CONNECT: eq50 0 0 0 0 @eq 0 0 1 50
// Retrieval info: CONNECT: eq51 0 0 0 0 @eq 0 0 1 51
// Retrieval info: CONNECT: eq52 0 0 0 0 @eq 0 0 1 52
// Retrieval info: CONNECT: eq53 0 0 0 0 @eq 0 0 1 53
// Retrieval info: CONNECT: eq54 0 0 0 0 @eq 0 0 1 54
// Retrieval info: CONNECT: eq55 0 0 0 0 @eq 0 0 1 55
// Retrieval info: CONNECT: eq56 0 0 0 0 @eq 0 0 1 56
// Retrieval info: CONNECT: eq57 0 0 0 0 @eq 0 0 1 57
// Retrieval info: CONNECT: eq58 0 0 0 0 @eq 0 0 1 58
// Retrieval info: CONNECT: eq59 0 0 0 0 @eq 0 0 1 59
// Retrieval info: CONNECT: eq6 0 0 0 0 @eq 0 0 1 6
// Retrieval info: CONNECT: eq60 0 0 0 0 @eq 0 0 1 60
// Retrieval info: CONNECT: eq61 0 0 0 0 @eq 0 0 1 61
// Retrieval info: CONNECT: eq62 0 0 0 0 @eq 0 0 1 62
// Retrieval info: CONNECT: eq63 0 0 0 0 @eq 0 0 1 63
// Retrieval info: CONNECT: eq7 0 0 0 0 @eq 0 0 1 7
// Retrieval info: CONNECT: eq8 0 0 0 0 @eq 0 0 1 8
// Retrieval info: CONNECT: eq9 0 0 0 0 @eq 0 0 1 9
// Retrieval info: GEN_FILE: TYPE_NORMAL peripheral_addr_dec.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL peripheral_addr_dec.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL peripheral_addr_dec.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL peripheral_addr_dec.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL peripheral_addr_dec_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL peripheral_addr_dec_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
